netcdf testrh {
dimensions:
	dim1 = 10000 ;
variables:
	float var1(dim1) ;
data:

 var1 = 420, 197, 391.5, 399, 455.5, 98.5, 167.5, 384, 138.5, 276.5, 238.5, 
    314, 182, 256.5, 476, 458, 317.5, 358.5, 70.5, 303, 8, 121, 68.5, 402, 
    78, 200, 64.5, 54, 499, 109, 256, 419.5, 306, 148, 318.5, 262, 246.5, 
    486, 146, 385.5, 263, 384.5, 200, 445.5, 141.5, 176, 403.5, 459.5, 34.5, 
    474.5, 262.5, 43, 96, 331.5, 445, 174, 32, 10, 228.5, 31.5, 119, 485, 
    451, 425, 133, 269.5, 187.5, 380, 256, 333.5, 265.5, 19.5, 218.5, 465.5, 
    465, 360, 142, 369, 319.5, 177, 343.5, 82.5, 220, 440, 414.5, 165, 114, 
    446.5, 175, 343, 478, 294, 328.5, 429, 219.5, 461.5, 199, 407, 342, 455, 
    241, 107.5, 475, 460, 73.5, 440.5, 320.5, 215.5, 309.5, 140.5, 393, 
    153.5, 223.5, 113, 93.5, 138, 278, 208, 84.5, 453, 51.5, 63, 247.5, 380, 
    492, 467.5, 342, 191.5, 374.5, 184, 147, 116, 292, 122, 76, 366, 62.5, 
    396.5, 82, 372.5, 37, 475, 26, 260.5, 88, 120, 398.5, 366, 328, 483.5, 
    319.5, 379.5, 46.5, 67, 260, 39, 34.5, 102, 230.5, 409.5, 286.5, 377.5, 
    25.5, 78.5, 499.5, 102, 444.5, 62.5, 498.5, 27, 435, 36, 2, 461.5, 296.5, 
    90, 81.5, 195.5, 456.5, 409.5, 179.5, 276, 289.5, 226, 343.5, 49.5, 265, 
    378.5, 152, 496, 288, 438.5, 373.5, 314, 17.5, 373.5, 416.5, 462.5, 
    436.5, 415.5, 489.5, 371.5, 451.5, 491.5, 333, 248.5, 81.5, 415, 444, 38, 
    324.5, 124, 314.5, 114.5, 350, 158, 164, 115.5, 37, 316.5, 111.5, 325.5, 
    255, 485.5, 140, 273, 359.5, 56.5, 235.5, 296, 472, 225, 168, 423.5, 217, 
    1.5, 172, 299, 416.5, 116.5, 337.5, 241, 240.5, 152, 356, 91, 310.5, 20, 
    206.5, 347.5, 336.5, 318.5, 173.5, 92, 304.5, 313.5, 365, 164, 370, 101, 
    460, 342, 326.5, 128.5, 266, 43.5, 130, 438.5, 343, 46.5, 55.5, 180.5, 
    288, 296.5, 333, 144, 387.5, 144, 164.5, 94.5, 492, 1.5, 413.5, 165.5, 
    94, 218, 479, 459, 382, 349.5, 60.5, 342.5, 191.5, 387, 471.5, 458, 
    430.5, 101.5, 396.5, 274, 148.5, 452, 454.5, 436.5, 249, 288, 81, 136.5, 
    432, 246, 231.5, 424, 247.5, 145.5, 90, 342, 363.5, 69.5, 301.5, 246, 
    419, 362, 89, 110.5, 249, 60.5, 69, 180, 162, 465.5, 454, 311, 418, 409, 
    248, 167, 197, 329, 304, 129, 75.5, 36, 53.5, 323.5, 181.5, 144, 165.5, 
    45.5, 213.5, 467, 291.5, 132.5, 329, 380.5, 243.5, 78.5, 441.5, 312.5, 
    258.5, 103.5, 278.5, 213, 414.5, 197, 122, 163, 364.5, 319, 492, 169, 
    448.5, 68, 205, 2.5, 391.5, 387, 146.5, 57, 432.5, 360.5, 24.5, 224.5, 
    493, 353.5, 105, 236.5, 432.5, 46.5, 49.5, 191, 150.5, 328.5, 404.5, 
    65.5, 25.5, 26.5, 228.5, 390, 346, 221, 59.5, 294.5, 289, 264.5, 297.5, 
    180.5, 152, 444, 238, 84.5, 304.5, 262.5, 309, 298, 116.5, 414.5, 35, 49, 
    461.5, 84.5, 240.5, 112.5, 413, 145, 178.5, 439, 172, 407, 329.5, 18, 
    128.5, 389, 312.5, 418, 154, 110.5, 99, 306, 54.5, 337, 391, 359.5, 100, 
    200.5, 157.5, 217, 115, 192.5, 266, 77, 277.5, 7, 190, 191, 152.5, 368.5, 
    130, 324.5, 276, 459.5, 342.5, 404.5, 348.5, 155.5, 322.5, 3, 266, 421.5, 
    309, 321, 259, 200, 181, 359, 400.5, 338.5, 76, 16, 31.5, 342.5, 93.5, 
    309, 350, 283.5, 0.5, 2.5, 152.5, 130.5, 327.5, 428.5, 90.5, 170.5, 
    333.5, 439.5, 326.5, 156.5, 442.5, 93, 78.5, 251.5, 414, 337.5, 452, 
    95.5, 197, 353, 434, 273.5, 369, 466, 116.5, 463, 275.5, 466.5, 247, 276, 
    469.5, 399.5, 407, 297, 328.5, 497.5, 467.5, 162, 437, 294.5, 318.5, 
    379.5, 387.5, 397, 131, 302, 235, 83, 397.5, 432.5, 436.5, 332, 206, 
    305.5, 298, 322.5, 269, 74, 289.5, 16, 350, 259, 416, 257.5, 56, 244.5, 
    255, 24, 407, 192, 318.5, 226, 71.5, 206.5, 123.5, 203, 8.5, 358.5, 
    286.5, 406, 291, 223, 238.5, 497.5, 29, 37, 320, 298.5, 111, 109.5, 315, 
    461.5, 368.5, 231, 219, 425, 476, 474, 449.5, 383.5, 166.5, 268, 109.5, 
    238.5, 474.5, 233, 442, 483.5, 91.5, 229, 390, 383, 452, 128.5, 380.5, 
    481.5, 165.5, 201, 280, 277, 311, 95.5, 238.5, 180, 326.5, 458, 105, 303, 
    432.5, 54.5, 186.5, 99.5, 323, 296, 338, 298, 29, 280, 281.5, 121, 9, 
    171.5, 4.5, 461.5, 300.5, 385, 443.5, 466.5, 86.5, 223.5, 243.5, 397.5, 
    319.5, 482.5, 77.5, 146, 441, 183, 449.5, 373.5, 237.5, 136, 473, 61, 
    432.5, 311.5, 359, 462, 92, 141, 83.5, 101, 313, 88, 63, 113.5, 473, 6.5, 
    80, 59.5, 230.5, 324, 457.5, 50, 307, 35, 196.5, 248, 218, 146.5, 122, 
    456, 283, 95, 17, 215.5, 406.5, 376.5, 178, 498.5, 17.5, 261.5, 100, 
    330.5, 349.5, 163.5, 444.5, 323, 170.5, 25, 383, 401.5, 349, 340.5, 452, 
    156, 376, 148.5, 404.5, 94.5, 295.5, 26.5, 50.5, 78.5, 122, 68, 294.5, 
    29, 444.5, 472.5, 28, 462.5, 234.5, 128, 293.5, 84, 292, 238, 407.5, 463, 
    263, 291, 364.5, 112.5, 132, 316.5, 269, 8, 465.5, 173.5, 102.5, 261, 
    200, 153.5, 339.5, 322.5, 221.5, 134.5, 351.5, 166, 107, 379.5, 129, 
    341.5, 8, 422.5, 426, 300, 160.5, 333.5, 263, 424, 125, 128, 36.5, 257, 
    444.5, 305.5, 265.5, 410.5, 479, 368, 171.5, 179.5, 21.5, 11.5, 2.5, 
    243.5, 146, 354, 410, 253.5, 233.5, 39, 95, 241.5, 461.5, 21.5, 42, 122, 
    355.5, 305.5, 46, 480.5, 433.5, 83, 237.5, 378.5, 388.5, 3, 289, 368, 
    371.5, 461, 48, 393.5, 473, 50.5, 137, 119.5, 404.5, 47.5, 373, 138.5, 
    86.5, 468.5, 380, 48, 490.5, 422.5, 170.5, 346, 228, 217, 327, 161.5, 
    300, 64.5, 40.5, 188.5, 68, 329.5, 57, 440, 291, 105, 334, 264, 156, 
    471.5, 384, 61, 19, 257, 199.5, 105.5, 226, 80, 154, 216.5, 2.5, 324.5, 
    63, 230.5, 42, 390, 392.5, 342, 455, 433.5, 31, 23.5, 263.5, 88.5, 463.5, 
    54.5, 193.5, 298, 319, 350, 269.5, 203, 411, 288.5, 460.5, 110.5, 394.5, 
    187, 190.5, 48.5, 403.5, 193.5, 373.5, 467, 424.5, 415.5, 357, 317.5, 
    258, 312, 251, 289, 335.5, 14.5, 377.5, 299.5, 69.5, 71.5, 97.5, 388.5, 
    422, 367.5, 92, 333, 156, 52.5, 444, 51, 239.5, 135, 99.5, 143.5, 328.5, 
    473.5, 110.5, 253, 389, 468, 71, 147, 280.5, 322, 436.5, 116, 336.5, 
    314.5, 416, 406, 386.5, 14, 295, 308.5, 381.5, 387, 142, 38, 440, 86, 89, 
    179.5, 221.5, 189, 323.5, 50, 162.5, 434.5, 303.5, 52, 402.5, 374.5, 199, 
    183, 197, 136, 299.5, 34, 450.5, 216, 440.5, 337, 230, 235.5, 146, 112, 
    123, 288, 150.5, 63, 374.5, 240, 242.5, 96, 429, 66.5, 146.5, 92, 1, 450, 
    144, 404, 325, 343.5, 87.5, 22, 479.5, 387.5, 56, 430.5, 103.5, 497, 268, 
    333.5, 232.5, 414, 446, 355.5, 202.5, 96.5, 418.5, 77, 336.5, 161.5, 
    173.5, 266, 228.5, 320, 358.5, 230, 270.5, 2.5, 134, 95.5, 346.5, 222, 
    118, 326.5, 109.5, 174.5, 257, 213, 171.5, 25, 47, 404.5, 439.5, 493, 
    260.5, 142, 90, 179.5, 219, 426.5, 341.5, 393, 193, 70, 213, 51.5, 300, 
    483.5, 54.5, 434.5, 79.5, 401, 156.5, 197.5, 227.5, 266, 372.5, 485, 479, 
    44, 10, 26.5, 448.5, 449.5, 19.5, 209.5, 91.5, 109.5, 389, 311, 36.5, 
    230.5, 204, 229.5, 300.5, 417.5, 281.5, 101, 401.5, 336, 35.5, 481, 
    237.5, 192, 179, 465, 458, 51.5, 450, 437.5, 95.5, 460.5, 464, 44.5, 410, 
    484, 254, 2, 94, 143.5, 313.5, 130.5, 374, 18, 360.5, 175, 436, 142.5, 
    276, 337.5, 478.5, 312, 318.5, 216, 4, 498, 181.5, 462.5, 49.5, 132, 
    400.5, 145.5, 93, 364.5, 190, 3, 349, 444.5, 5.5, 443, 88, 319.5, 74, 
    462.5, 337.5, 435, 137.5, 273.5, 77.5, 414, 111, 56, 226, 430, 272.5, 
    230.5, 428, 454.5, 193, 478, 87, 93.5, 123.5, 180, 458.5, 313.5, 183.5, 
    307.5, 258.5, 189, 250.5, 347, 8.5, 325, 309.5, 346.5, 260, 447.5, 120.5, 
    337.5, 361.5, 232, 394, 88, 162.5, 167, 318.5, 91, 121.5, 12, 69, 208.5, 
    106, 192.5, 388.5, 64.5, 6.5, 72, 372.5, 265, 261.5, 123, 112, 270.5, 
    448.5, 422, 117.5, 208.5, 369.5, 238, 46, 231.5, 470.5, 440, 320, 133, 
    107, 139, 224, 229, 151, 293, 437.5, 257, 485.5, 326.5, 322, 492, 399, 
    194.5, 257.5, 161, 318, 370, 432, 266.5, 292, 49.5, 475, 161.5, 288, 
    21.5, 393.5, 258.5, 462, 213.5, 392, 69, 352.5, 116, 298.5, 3.5, 409.5, 
    236.5, 261, 395, 63, 83.5, 387.5, 462.5, 278, 145.5, 123.5, 96.5, 15.5, 
    56, 363.5, 307.5, 105.5, 339, 469.5, 394, 360.5, 363, 152.5, 322.5, 77, 
    45, 392, 429.5, 161, 190.5, 433.5, 70.5, 427, 195, 466, 490.5, 278.5, 
    354, 453, 57, 0, 77, 153.5, 15.5, 133.5, 17.5, 323.5, 239, 356.5, 293.5, 
    133.5, 217, 157, 286.5, 40, 234, 331.5, 432, 163.5, 492.5, 123, 97, 63.5, 
    50.5, 292, 30, 41, 71, 384.5, 494.5, 128, 384.5, 72, 282, 400, 205.5, 
    299.5, 224, 445, 156, 17.5, 78.5, 373.5, 174.5, 365, 413.5, 408.5, 196.5, 
    346, 72.5, 189.5, 469, 170, 253.5, 20, 462.5, 284, 61, 33.5, 168.5, 56, 
    162, 53, 128, 444, 453.5, 334, 243.5, 177.5, 279, 400, 195, 358, 273.5, 
    370, 223, 187, 279, 420, 33.5, 351.5, 110, 3, 21.5, 364, 23, 484.5, 148, 
    84.5, 18, 316.5, 140.5, 180, 369.5, 269, 124.5, 323, 103, 368, 1, 382, 
    268.5, 196.5, 240.5, 42, 66.5, 464, 229.5, 345.5, 384, 263, 197.5, 494.5, 
    266.5, 219.5, 358.5, 289.5, 204, 7, 374, 222.5, 323.5, 15, 403, 193.5, 
    284, 27.5, 17, 387, 396, 18, 269.5, 164.5, 214.5, 10, 206.5, 281.5, 474, 
    436.5, 127, 358.5, 199.5, 325, 353, 466.5, 44.5, 212, 256, 248.5, 219, 
    130.5, 471.5, 43, 146, 374.5, 237, 430, 402, 254, 317.5, 298, 272, 87, 
    463, 487, 97.5, 170, 268.5, 72, 106.5, 396, 430.5, 306.5, 221, 284, 273, 
    266, 496.5, 29.5, 15, 216, 160.5, 486.5, 259.5, 306.5, 361, 496.5, 236.5, 
    263.5, 250.5, 54.5, 61.5, 23, 141.5, 25, 10, 239.5, 195, 279, 311.5, 
    301.5, 175.5, 242.5, 108, 396.5, 27, 381, 163, 23.5, 410.5, 178, 240, 71, 
    164.5, 499.5, 378, 25.5, 496, 114.5, 289, 246.5, 169.5, 351, 270, 311, 
    376, 280.5, 51, 71.5, 59.5, 363, 373, 235, 105.5, 481.5, 132, 132.5, 
    362.5, 295, 156.5, 273.5, 473, 396.5, 345, 138, 396, 223, 163.5, 392.5, 
    338, 453, 139.5, 7.5, 304.5, 409.5, 319, 181, 190, 370.5, 252.5, 250, 
    233.5, 125.5, 485, 339, 107.5, 117.5, 472, 470, 412.5, 129, 244, 386, 26, 
    89, 24, 422.5, 312.5, 188, 315, 151, 141.5, 454.5, 158.5, 446, 364, 478, 
    127, 54.5, 348.5, 379.5, 304.5, 82.5, 5.5, 290, 421.5, 113, 407.5, 394, 
    83.5, 320.5, 23, 328, 206.5, 49, 417.5, 231, 471.5, 230, 419.5, 287, 381, 
    61, 241.5, 40, 7, 106, 18.5, 134.5, 160.5, 367.5, 14.5, 465.5, 450, 20, 
    255.5, 372, 133.5, 163, 266, 217.5, 483.5, 289.5, 45.5, 190.5, 339, 463, 
    422, 311, 193.5, 341.5, 98, 74.5, 403, 340, 115, 410.5, 446, 134, 45, 
    107, 1.5, 59.5, 73, 451.5, 80, 328.5, 323.5, 213.5, 492, 90, 431, 476, 
    379.5, 477, 166.5, 218.5, 440, 89, 30, 133.5, 431, 128, 208.5, 334, 468, 
    324, 244.5, 414.5, 458, 289.5, 22, 459.5, 349.5, 95, 411, 429.5, 424, 
    235, 143.5, 416, 325, 75, 392, 205, 52, 59, 423.5, 492, 148, 454, 126, 
    79, 82, 335, 413.5, 50.5, 159, 158, 465.5, 117, 448, 487.5, 76.5, 297.5, 
    82.5, 488, 227.5, 6.5, 223.5, 371, 423, 48.5, 446, 315, 253.5, 498.5, 
    374, 177.5, 490.5, 22, 131.5, 117, 101.5, 214, 452, 15, 264.5, 111, 
    173.5, 230, 228.5, 121.5, 218, 305.5, 419.5, 301, 293.5, 147.5, 307.5, 
    17.5, 18.5, 231, 66, 465, 46, 320, 463.5, 420.5, 497.5, 454.5, 443, 
    129.5, 72, 44.5, 343.5, 24, 60, 108.5, 135.5, 233.5, 339, 364, 355.5, 57, 
    169.5, 275.5, 358, 463.5, 423, 166, 481, 442, 397, 47.5, 407.5, 443, 
    367.5, 371, 363.5, 365, 326, 306.5, 495, 398, 351.5, 338.5, 422.5, 411.5, 
    447.5, 58, 145.5, 286.5, 422.5, 1, 343.5, 92.5, 276.5, 201.5, 56, 200, 
    367.5, 37.5, 142.5, 264.5, 85, 50, 208, 453, 421.5, 72, 318.5, 247.5, 
    379, 313.5, 146, 230.5, 152, 69, 142.5, 99.5, 127.5, 288, 386.5, 50, 
    289.5, 230, 143, 66.5, 431.5, 199.5, 266.5, 299.5, 237, 409, 64.5, 322.5, 
    459, 273, 275.5, 381, 345, 94, 128.5, 224.5, 407.5, 275, 455, 60, 344, 
    98, 160, 471.5, 386, 46.5, 22, 175.5, 277, 165, 242, 208.5, 364.5, 9, 
    8.5, 102, 418.5, 73.5, 424.5, 378, 346.5, 200.5, 259, 192, 295, 388, 
    416.5, 202.5, 163, 371.5, 263, 7.5, 469.5, 423.5, 479.5, 356, 470.5, 1.5, 
    32, 247.5, 166.5, 274.5, 456.5, 31.5, 283.5, 465, 133.5, 202.5, 38.5, 
    58.5, 80.5, 385.5, 259, 339.5, 77.5, 54, 228, 494, 257, 391.5, 366, 20.5, 
    399, 336, 444, 378.5, 192, 415, 380.5, 224, 162.5, 47, 499, 119, 79, 
    282.5, 84.5, 212.5, 485.5, 123.5, 271.5, 66, 9, 30.5, 406, 87, 85, 134, 
    81, 342, 25.5, 447, 363, 424.5, 283, 307, 303.5, 475.5, 222.5, 184, 200, 
    385, 231.5, 199, 4.5, 310.5, 482, 89.5, 23.5, 467.5, 213, 295, 33.5, 
    222.5, 326, 439.5, 310, 411, 74, 391, 253.5, 99.5, 338.5, 116.5, 24.5, 
    122, 424, 328, 97.5, 146.5, 12.5, 297.5, 32, 244, 496.5, 37, 55, 479, 
    126.5, 79, 446.5, 340, 374, 480.5, 63, 200.5, 420, 373, 112, 494.5, 264, 
    365.5, 94, 103, 482.5, 119, 225, 407, 447.5, 322.5, 54, 460, 120, 86.5, 
    204.5, 117, 123.5, 259.5, 96, 250, 338.5, 43, 90, 213, 23.5, 153, 413.5, 
    443.5, 26, 25.5, 438.5, 290.5, 391.5, 32.5, 393.5, 374.5, 152, 118.5, 
    282, 99.5, 441.5, 336.5, 59.5, 62, 423, 264, 179, 47, 24, 275.5, 297, 
    363, 318.5, 387.5, 76, 342, 41, 490, 286, 67.5, 16, 224.5, 358.5, 407.5, 
    257.5, 252, 282.5, 409.5, 371, 65, 9, 313, 401.5, 69, 375, 325, 333.5, 
    54.5, 372, 358, 330, 169, 221, 149, 57, 297, 491.5, 98.5, 287.5, 278, 
    166, 303.5, 3, 24.5, 211.5, 260.5, 277, 494.5, 170.5, 148.5, 59.5, 180, 
    461.5, 461, 249.5, 337, 286, 83, 391.5, 158, 441, 222, 327.5, 162.5, 
    371.5, 385, 460, 363, 483.5, 247.5, 141, 150, 51, 144, 175, 263, 405, 
    452.5, 257.5, 76, 101, 317, 256.5, 63, 278.5, 6, 400, 64.5, 89.5, 292, 
    223, 31, 14, 51, 193.5, 385.5, 436, 153.5, 249, 420, 401, 390, 70, 452.5, 
    34.5, 245, 215.5, 440, 197.5, 473, 16.5, 299, 290, 273, 362.5, 68.5, 279, 
    263, 133.5, 368.5, 55, 357, 399.5, 69, 408, 93, 455, 344.5, 247, 204, 
    264.5, 148, 94.5, 335, 101, 129.5, 80.5, 316.5, 70, 278.5, 290, 86.5, 78, 
    80.5, 359.5, 440.5, 149.5, 138.5, 203.5, 283, 7.5, 258.5, 140, 407.5, 
    328, 48.5, 1, 283, 393.5, 248, 487.5, 158, 396.5, 82, 493.5, 497.5, 
    211.5, 74.5, 314.5, 282, 353, 104.5, 368.5, 431, 185, 228, 372, 334.5, 
    367, 76, 118, 375, 334.5, 258.5, 282.5, 163, 307, 283.5, 446.5, 200.5, 
    31.5, 434, 359, 428.5, 16.5, 353, 426, 228.5, 427.5, 241, 10.5, 280.5, 
    346, 379, 212, 31, 107.5, 84.5, 366, 474.5, 160.5, 484.5, 349.5, 495.5, 
    243, 132, 158.5, 50.5, 416, 105, 251.5, 447.5, 39.5, 111, 376, 56, 464, 
    302.5, 284.5, 392, 44, 295, 172.5, 390, 174, 385, 421.5, 281.5, 469.5, 
    288, 256.5, 130, 272.5, 106.5, 126, 16, 238.5, 284.5, 66.5, 154.5, 390, 
    318, 102.5, 429.5, 429.5, 479, 486, 393.5, 282, 270.5, 285.5, 326, 65.5, 
    458.5, 216.5, 240, 344, 138, 22, 314, 426, 279, 444.5, 198.5, 385.5, 
    70.5, 214.5, 124.5, 355, 281.5, 279.5, 245.5, 100, 382.5, 175, 29.5, 
    361.5, 161, 423.5, 144, 432, 209, 470.5, 498, 168, 187, 238.5, 12, 325, 
    261, 326.5, 251.5, 40, 271, 450, 425.5, 341.5, 165, 50.5, 197, 446.5, 
    330, 442.5, 47, 212.5, 118, 76.5, 74.5, 279.5, 0, 218.5, 211.5, 209.5, 
    189, 210, 377.5, 376.5, 448.5, 390, 202, 209.5, 216.5, 453.5, 250, 487.5, 
    404, 175.5, 329.5, 69, 226, 26.5, 16, 56.5, 469.5, 63, 269, 87.5, 140, 
    343.5, 367, 140, 62.5, 79, 349.5, 252, 289, 227.5, 128.5, 238, 118, 
    330.5, 448, 334.5, 284.5, 198, 322.5, 188.5, 373.5, 152.5, 258, 100, 179, 
    274, 157, 148.5, 337.5, 426, 236.5, 477.5, 270, 104, 118, 332.5, 183, 
    468, 85, 472.5, 195.5, 213.5, 210.5, 313.5, 44.5, 159, 148.5, 329.5, 357, 
    471.5, 18, 231, 124, 276, 331, 303.5, 50.5, 488, 452, 388.5, 414.5, 189, 
    366.5, 184.5, 293, 484.5, 17.5, 476.5, 453, 102.5, 449, 148.5, 316.5, 
    160, 462.5, 361.5, 319, 111.5, 191.5, 176, 83, 209.5, 407, 207.5, 486, 
    238.5, 11, 36.5, 227, 463.5, 425.5, 142, 152.5, 292, 327, 446, 277, 345, 
    422.5, 230, 448, 372, 379, 265, 32.5, 342, 126.5, 351.5, 453.5, 318, 28, 
    37, 28, 435.5, 244.5, 14, 174.5, 255.5, 51, 402, 219.5, 476.5, 44, 372, 
    269, 371.5, 318, 46, 216.5, 241, 276.5, 164.5, 113, 155.5, 429.5, 145.5, 
    497.5, 56.5, 497.5, 451.5, 375, 26, 489, 403, 462, 233.5, 417.5, 136.5, 
    489.5, 468.5, 39, 209, 445.5, 83.5, 81.5, 214.5, 455, 400, 261, 171.5, 
    141, 37.5, 336, 254, 193.5, 266, 400, 191, 322.5, 397.5, 143, 197.5, 
    423.5, 132, 101, 385.5, 366, 18.5, 22.5, 356, 487.5, 61.5, 65.5, 433, 
    145, 147, 148, 100.5, 47.5, 409, 272, 188.5, 447, 108.5, 443, 140.5, 
    374.5, 343, 332, 197, 241, 475, 395, 165, 107.5, 496, 50.5, 474, 15, 
    73.5, 330, 2.5, 135.5, 395.5, 436, 280.5, 43, 84.5, 381, 91, 494, 153.5, 
    279.5, 441.5, 262, 223, 82, 137, 66.5, 414, 334.5, 308, 389.5, 229.5, 
    473, 497.5, 226, 24, 471.5, 241, 97.5, 301.5, 244, 233, 197.5, 180.5, 14, 
    241, 265.5, 395.5, 332, 259.5, 49.5, 112, 201, 312, 335, 283.5, 449, 402, 
    197.5, 283.5, 210, 87.5, 13.5, 183.5, 85, 239.5, 207.5, 57, 481, 305.5, 
    359, 225.5, 39, 57, 406, 53, 298, 172, 449, 130, 432, 498.5, 242.5, 133, 
    311, 78, 417, 260, 480, 115, 44, 190.5, 202.5, 57.5, 374, 288, 297.5, 82, 
    345, 278.5, 387.5, 204.5, 4, 426.5, 261.5, 410.5, 480, 59.5, 82.5, 429.5, 
    190, 14.5, 428.5, 432.5, 148, 239.5, 11, 65, 499.5, 491.5, 180.5, 43.5, 
    182, 383, 101.5, 56.5, 171.5, 399, 138.5, 17, 177.5, 26.5, 221.5, 182, 
    453.5, 483, 93, 433.5, 43, 176, 363.5, 233.5, 191, 292, 166.5, 339.5, 
    31.5, 177.5, 405, 31.5, 169, 85.5, 75.5, 351.5, 469, 177, 408, 140.5, 76, 
    47, 158, 254, 74, 379.5, 436.5, 27.5, 363, 29.5, 461.5, 406.5, 206, 325, 
    140, 397, 117.5, 306.5, 237, 149, 484.5, 142, 180.5, 153.5, 227.5, 256, 
    5, 196.5, 433.5, 413.5, 337.5, 9.5, 460.5, 495.5, 264, 34.5, 375.5, 
    200.5, 62.5, 238.5, 230.5, 24, 145.5, 436.5, 349.5, 285.5, 334, 467, 
    92.5, 71, 116, 77, 213, 297, 230.5, 441, 53.5, 236, 138, 487, 149.5, 
    475.5, 497, 110.5, 471.5, 261, 145.5, 347.5, 461.5, 208, 86.5, 192.5, 
    232.5, 232, 129, 82, 17.5, 463, 49, 110.5, 34, 165.5, 187.5, 247.5, 463, 
    418.5, 188.5, 17, 154.5, 326.5, 4.5, 304.5, 302.5, 1.5, 415.5, 274.5, 
    263, 61, 122, 225, 269.5, 208.5, 417.5, 2, 440.5, 46.5, 84.5, 458.5, 10, 
    134, 69, 44.5, 300, 257, 292, 263.5, 175.5, 481, 280.5, 330.5, 307.5, 
    285.5, 135.5, 110.5, 287, 51, 385, 50.5, 112.5, 7.5, 275.5, 382, 216, 
    193.5, 384.5, 156.5, 240, 469.5, 115.5, 250.5, 104, 184.5, 295, 404, 
    441.5, 87, 167.5, 117.5, 68, 448.5, 448, 376, 234, 84, 487, 21.5, 135, 
    372.5, 72, 248, 380, 348, 130.5, 96, 41.5, 15, 253, 282, 485, 368.5, 
    32.5, 89, 53.5, 327.5, 493, 495.5, 415, 161, 113, 483.5, 110, 61.5, 360, 
    344, 146, 347, 365.5, 281, 220, 438, 29.5, 100, 286.5, 160, 196, 328, 
    175.5, 449.5, 110.5, 160.5, 318.5, 143, 249.5, 372, 471, 243, 368, 386.5, 
    404.5, 481, 370.5, 14.5, 43, 230.5, 359, 189, 78, 225, 470.5, 298, 163, 
    0, 398.5, 450, 160, 95, 278, 336, 44.5, 389, 496.5, 363, 32, 246.5, 
    235.5, 3.5, 490, 103.5, 390.5, 394.5, 85, 261, 409.5, 128.5, 492, 268.5, 
    318, 70.5, 493.5, 289, 369, 157, 289, 267.5, 107, 449.5, 362.5, 385.5, 
    285.5, 407.5, 274.5, 282.5, 271, 307, 29, 6.5, 311, 19.5, 110.5, 201.5, 
    414.5, 196, 462.5, 324, 324.5, 455, 92.5, 142.5, 25.5, 86.5, 431.5, 
    394.5, 243.5, 221, 162, 351, 171, 25, 236.5, 457, 432.5, 11.5, 239.5, 
    203.5, 318.5, 269, 210.5, 130, 288.5, 321.5, 331.5, 203, 17.5, 294.5, 27, 
    342.5, 249.5, 120, 485.5, 275, 207, 417, 169.5, 451, 138.5, 332, 302, 
    309.5, 357, 39, 267, 290, 50.5, 6.5, 494, 369.5, 275.5, 205, 499.5, 64, 
    26.5, 331.5, 267, 44.5, 126, 294.5, 387, 375.5, 415, 372.5, 151, 122, 
    290, 321, 73, 428.5, 153.5, 375.5, 238.5, 10.5, 414.5, 5.5, 301, 465.5, 
    12.5, 295, 335.5, 288, 0, 335, 352.5, 27, 166.5, 120, 71.5, 293, 414.5, 
    458.5, 169, 329.5, 331.5, 320, 452, 121.5, 141.5, 25, 50.5, 295, 401, 
    289.5, 306, 316, 295.5, 107, 281.5, 308, 402, 117, 96.5, 402.5, 452.5, 
    449.5, 430, 119.5, 69.5, 1.5, 412.5, 484, 460.5, 81.5, 314, 292.5, 402, 
    266.5, 414, 43.5, 292, 465, 339, 193, 255, 145, 9, 51, 252, 290.5, 359.5, 
    154.5, 408, 456, 57.5, 361, 405.5, 487.5, 480.5, 475, 489.5, 393.5, 
    459.5, 450.5, 475, 274, 243, 377.5, 40.5, 157.5, 421.5, 333, 123, 260.5, 
    26, 378, 406, 35, 429, 158, 326, 288.5, 313, 234.5, 245, 371, 95.5, 151, 
    358.5, 76, 126.5, 348.5, 469.5, 86.5, 299.5, 445, 360.5, 42.5, 323, 
    401.5, 200.5, 244.5, 234.5, 324, 5.5, 261, 202, 411.5, 296, 131.5, 69.5, 
    122.5, 420.5, 383, 357.5, 166, 254, 453, 317, 113, 29.5, 443.5, 462, 
    499.5, 30, 261.5, 445, 391, 304.5, 268, 293, 5, 12.5, 27.5, 329, 18, 289, 
    31.5, 429.5, 85, 163.5, 499.5, 208, 84, 382.5, 65.5, 250.5, 137, 19, 
    67.5, 250, 48.5, 11.5, 212, 48.5, 42, 474, 493.5, 433, 278.5, 261.5, 
    226.5, 283.5, 274.5, 254.5, 113, 292.5, 43.5, 145, 222.5, 129, 308.5, 
    222.5, 337, 393, 105, 403, 143.5, 242.5, 422, 211.5, 493, 471, 223, 
    205.5, 19.5, 265, 179.5, 13, 198.5, 458, 275, 425.5, 242, 49.5, 180, 
    355.5, 342.5, 223.5, 0.5, 65, 352.5, 309, 287.5, 190, 202.5, 393, 93, 
    346, 136, 15.5, 57.5, 129, 487, 281, 334.5, 6.5, 46.5, 14.5, 20, 245.5, 
    472.5, 295, 171, 215, 345, 351, 70.5, 187.5, 75, 71, 253, 427.5, 380.5, 
    41, 118, 83, 434, 211.5, 429.5, 70.5, 227.5, 487, 199.5, 214.5, 268.5, 
    34.5, 221, 315, 49, 241.5, 61, 21.5, 36.5, 232, 237, 381.5, 83, 307.5, 
    69.5, 158.5, 379, 322.5, 86.5, 260, 363.5, 204.5, 343.5, 298, 416.5, 273, 
    368.5, 144, 260.5, 68, 358.5, 29, 102.5, 80, 344.5, 152, 321.5, 405.5, 
    173.5, 358.5, 137.5, 411, 240, 221, 218.5, 310, 380, 98, 132.5, 466.5, 
    358.5, 496.5, 171, 202, 294.5, 88, 475, 163.5, 232, 236, 232, 91, 265, 
    335, 171, 110, 487, 492.5, 16, 161, 351, 153.5, 72, 91.5, 375, 291, 
    401.5, 255.5, 389, 34.5, 222, 247.5, 31, 393.5, 450, 325.5, 481.5, 425.5, 
    489.5, 214, 161.5, 221.5, 305, 426.5, 56.5, 476, 37, 43.5, 468.5, 53, 
    204.5, 320, 207, 276.5, 412, 82.5, 67.5, 313.5, 338, 457, 348, 60, 205, 
    379, 454, 155, 205, 435.5, 80.5, 194.5, 149.5, 242.5, 416.5, 454.5, 
    169.5, 473, 431, 206.5, 17, 399.5, 260, 221.5, 220, 467, 498.5, 132, 
    49.5, 66.5, 446, 388, 24, 294, 448.5, 229, 173.5, 402.5, 384.5, 379, 338, 
    465.5, 74, 488, 208, 490.5, 443, 377.5, 464, 374, 84.5, 481, 274, 344.5, 
    202.5, 494, 311.5, 201.5, 126.5, 361.5, 268, 72.5, 249.5, 292, 366.5, 
    198, 21.5, 40.5, 100.5, 406, 420, 439, 372, 494, 427.5, 80, 485, 370.5, 
    458, 449, 244.5, 42.5, 430, 18.5, 387.5, 133, 12.5, 199, 334.5, 139, 61, 
    103, 211.5, 310.5, 395, 78.5, 9, 417, 119.5, 110, 323.5, 40, 49.5, 195.5, 
    34.5, 477, 276, 19.5, 347.5, 234.5, 469, 92, 277, 399.5, 111, 164.5, 
    32.5, 124, 364, 367.5, 263, 425, 471, 475, 236, 366.5, 54, 245.5, 283.5, 
    174, 356, 107, 214, 405.5, 302.5, 248.5, 382.5, 79, 268.5, 230.5, 313.5, 
    238, 323, 91, 137.5, 434, 256, 170.5, 58, 120, 38.5, 321.5, 45.5, 9.5, 
    297, 282, 376, 351.5, 27.5, 159.5, 25.5, 384, 267, 240, 289.5, 70, 489, 
    172.5, 149, 257.5, 403, 462.5, 495.5, 226.5, 53.5, 133.5, 160.5, 309.5, 
    304, 219, 430, 342.5, 40.5, 475.5, 352, 337.5, 257.5, 228.5, 189.5, 
    285.5, 388, 215, 169.5, 155.5, 455.5, 459.5, 225.5, 444.5, 132, 374.5, 
    202.5, 35.5, 337, 198, 262, 391, 332, 423, 201, 136, 142, 131, 479, 183, 
    106.5, 331.5, 21, 364.5, 60, 210.5, 150.5, 448.5, 426, 320.5, 104, 381.5, 
    280, 329.5, 326, 412, 204, 28.5, 448, 41.5, 227, 210.5, 433, 59, 134, 
    134, 195.5, 276, 265, 174.5, 459.5, 372, 6, 480.5, 237, 66.5, 191.5, 388, 
    15, 117.5, 208.5, 119, 499, 488.5, 448.5, 325, 401, 153, 354, 349, 195, 
    81, 59.5, 128, 140.5, 193.5, 262.5, 336.5, 470, 28, 11, 430, 400.5, 17.5, 
    411, 137.5, 84, 102.5, 25.5, 99, 220, 234, 218.5, 219.5, 223, 167.5, 45, 
    124, 321, 399, 473, 16, 480.5, 33, 144.5, 121.5, 227, 407, 458, 197.5, 
    435.5, 469.5, 127.5, 336, 487.5, 38.5, 473.5, 71.5, 141.5, 499.5, 171, 
    362, 234, 390, 81.5, 457, 57.5, 126.5, 81, 378.5, 26, 54.5, 395, 7, 88, 
    39.5, 128.5, 315, 447, 86.5, 13, 382.5, 56, 141, 218.5, 44, 179.5, 192.5, 
    115.5, 321.5, 192.5, 287, 183.5, 426.5, 177, 265.5, 384, 235, 392, 465.5, 
    113.5, 418.5, 20, 8.5, 425.5, 108, 48.5, 54, 423.5, 496, 141, 436.5, 
    378.5, 197.5, 77.5, 97.5, 241.5, 257.5, 290.5, 357.5, 79, 483, 145, 263, 
    410, 322, 28.5, 294, 57.5, 421, 259.5, 171, 339.5, 280, 180, 265.5, 388, 
    229, 319.5, 311.5, 225, 461, 248, 103.5, 159, 326, 201.5, 400.5, 83.5, 
    492, 258.5, 162.5, 475, 403.5, 426, 385.5, 225.5, 454.5, 180, 283, 375.5, 
    440, 454.5, 215.5, 220, 135, 481, 108, 364, 301, 420, 89, 262, 168.5, 
    193, 421, 494.5, 394.5, 322, 78, 386.5, 80.5, 241, 362, 484, 167, 247.5, 
    210, 121.5, 428, 493.5, 497.5, 368, 448, 213, 88, 83.5, 194, 196.5, 
    447.5, 495.5, 116.5, 36.5, 257.5, 285, 229.5, 179, 280, 124, 1.5, 358, 
    11, 82, 99, 373.5, 66.5, 266.5, 121.5, 276.5, 388.5, 49.5, 270.5, 386, 
    417.5, 219, 99, 5.5, 302.5, 293.5, 202, 250, 289, 319, 287, 47, 104.5, 
    17, 226.5, 384.5, 141.5, 228, 242.5, 152.5, 310.5, 342, 26, 377.5, 109, 
    148, 154, 497.5, 197.5, 424.5, 383.5, 115, 143.5, 483, 121, 446.5, 277, 
    323.5, 196.5, 66.5, 142.5, 484, 113.5, 247.5, 1, 340.5, 132, 142.5, 69, 
    375, 295.5, 380, 217.5, 322, 257.5, 326.5, 470, 412, 324, 167.5, 336.5, 
    208, 283, 480.5, 191, 404, 427, 468, 228, 124, 34.5, 371, 108, 148.5, 
    118.5, 109.5, 489.5, 250.5, 252, 59, 126, 48, 439, 343.5, 370, 196.5, 
    170, 340, 108.5, 494.5, 8, 445.5, 202.5, 291, 426.5, 393.5, 195.5, 354, 
    362, 423.5, 478.5, 397, 294.5, 87, 46, 413, 196.5, 36, 164, 449, 95, 290, 
    497, 34, 134, 367.5, 231, 304, 207.5, 340, 299, 215.5, 286, 1.5, 7, 
    212.5, 395.5, 202.5, 67, 258, 126, 45.5, 155, 421, 133, 201.5, 334.5, 
    329.5, 237.5, 498.5, 279, 332.5, 289, 276, 367, 423, 143.5, 98.5, 227.5, 
    351.5, 438.5, 26.5, 67.5, 224.5, 28, 74.5, 437.5, 424, 277.5, 4.5, 182, 
    404, 50.5, 337, 325, 184, 39, 159.5, 13.5, 277, 158.5, 293, 110, 447.5, 
    69.5, 477, 371, 213.5, 75.5, 99, 65, 14.5, 125.5, 133, 239.5, 154, 208, 
    177, 78, 485.5, 182, 260, 390, 233, 97.5, 215, 417, 137, 375, 431, 414, 
    34, 224, 24, 482, 293.5, 1.5, 353, 7, 77, 452, 72.5, 92, 78, 205.5, 
    331.5, 232, 413.5, 8.5, 310.5, 399.5, 191, 71, 289.5, 424, 169, 5, 341, 
    306, 380.5, 272, 220, 414.5, 496.5, 244.5, 396.5, 290, 246, 249.5, 297, 
    323.5, 202, 369.5, 415.5, 280, 75.5, 247, 12.5, 489, 256, 323.5, 389, 
    447, 394.5, 178.5, 371.5, 63.5, 184, 212.5, 370, 64.5, 485, 90, 479, 
    481.5, 334.5, 376, 272, 80.5, 125.5, 69, 404.5, 328, 439, 320, 108.5, 
    14.5, 67.5, 121, 4, 323.5, 445, 393, 271, 339.5, 72, 142.5, 403.5, 256, 
    355.5, 273.5, 321, 340.5, 363.5, 300.5, 322.5, 198.5, 176.5, 94.5, 279.5, 
    302.5, 164, 184, 130.5, 103.5, 4.5, 239, 118.5, 72, 360.5, 122.5, 395.5, 
    306, 16, 166.5, 145.5, 88, 309, 49, 344.5, 164.5, 322.5, 166, 5.5, 186.5, 
    466.5, 328.5, 385.5, 143, 423, 165.5, 445.5, 87.5, 349.5, 76.5, 191, 354, 
    316, 309.5, 426, 177, 432.5, 322, 483, 448.5, 489, 128.5, 37, 298, 178, 
    382, 463, 1, 48, 469, 187.5, 14.5, 297.5, 73.5, 158, 221, 239, 103.5, 
    309, 89, 180, 0, 443, 496.5, 310, 369.5, 173.5, 243, 192, 156.5, 191.5, 
    181, 285.5, 229, 479.5, 463.5, 111, 442.5, 465, 159.5, 412, 153, 174.5, 
    209.5, 226.5, 332.5, 431, 465.5, 436, 240, 54.5, 116.5, 240.5, 498, 113, 
    51, 368, 287, 294, 60, 443.5, 486, 241, 229.5, 215, 220.5, 193, 326.5, 
    163.5, 158.5, 486, 75.5, 311.5, 160.5, 285.5, 38, 493, 216.5, 3.5, 429.5, 
    457, 58.5, 46.5, 198, 57, 160, 249, 425, 447, 43, 485.5, 391, 29, 227, 
    120.5, 244.5, 447.5, 314, 71.5, 111.5, 472.5, 57.5, 187, 284, 218.5, 473, 
    322, 212, 190, 326, 142, 147, 385, 188.5, 345, 442, 349, 94.5, 367.5, 
    296.5, 137.5, 353, 187.5, 167, 80, 308.5, 412, 28, 123, 483.5, 139.5, 
    95.5, 41.5, 327, 380, 260, 300.5, 202.5, 472.5, 490.5, 29, 114.5, 138, 
    414.5, 303.5, 483.5, 356.5, 152.5, 78, 224.5, 449.5, 216, 78, 137.5, 
    383.5, 158, 446, 295.5, 186.5, 69, 279, 326.5, 165, 321, 154, 45.5, 81.5, 
    454.5, 248, 54, 445.5, 277.5, 169, 83.5, 192, 472.5, 67, 49, 125.5, 
    145.5, 273.5, 75, 361.5, 351.5, 212.5, 245, 10, 159, 40.5, 197, 228.5, 
    320, 23.5, 394, 141, 178, 439.5, 222.5, 133, 188, 277, 78.5, 465.5, 446, 
    162, 157.5, 419, 229.5, 207, 44.5, 375, 480.5, 120, 236.5, 332.5, 333, 
    482, 343, 492, 22.5, 40.5, 221, 343, 64.5, 115, 484.5, 242.5, 54.5, 
    207.5, 375.5, 243, 484.5, 454, 208.5, 431, 116.5, 366.5, 350, 346.5, 
    73.5, 395, 222, 54.5, 15, 459, 387, 348, 441, 230.5, 340.5, 464, 271, 62, 
    307.5, 335.5, 177, 292, 78.5, 232, 0, 454, 475, 485, 408.5, 184, 416, 
    25.5, 50.5, 266.5, 372.5, 124.5, 161.5, 94.5, 179, 176.5, 53.5, 66.5, 25, 
    495, 297, 366, 459.5, 68.5, 428, 267, 404.5, 105.5, 59.5, 483, 338, 59.5, 
    437.5, 313.5, 44.5, 346.5, 497.5, 461, 372, 48.5, 227.5, 244.5, 173, 389, 
    339.5, 352.5, 66, 393.5, 419, 91, 388.5, 216, 457.5, 348, 285, 385.5, 
    115, 189.5, 491.5, 175, 172.5, 329.5, 234.5, 110.5, 143, 279.5, 457, 141, 
    241, 329, 190, 468.5, 74, 363.5, 358, 413.5, 216, 424, 307, 135, 15.5, 
    196, 351.5, 473, 44, 136.5, 359, 159.5, 326.5, 351, 334.5, 499.5, 180.5, 
    69.5, 110, 324, 349, 67, 465.5, 90.5, 396, 155.5, 59, 470.5, 19.5, 417.5, 
    384, 235.5, 341.5, 191.5, 371, 357.5, 387.5, 222.5, 331, 432, 359.5, 190, 
    92, 186.5, 41, 427, 186, 222, 497, 296, 46.5, 346.5, 363, 12, 437, 259, 
    168, 496, 229.5, 187.5, 414, 114, 423.5, 255.5, 306, 294.5, 113.5, 194, 
    17.5, 444.5, 126, 377, 135, 218.5, 63.5, 176.5, 146, 249.5, 399, 143, 
    45.5, 445.5, 489.5, 409, 458, 426.5, 168, 126.5, 423, 398, 314, 337, 
    12.5, 238, 93, 318.5, 32.5, 206.5, 12.5, 50, 151.5, 139, 427.5, 286.5, 
    357.5, 491, 463.5, 3.5, 241, 362.5, 147, 287, 308.5, 136.5, 196, 266.5, 
    63, 364.5, 393, 486, 263, 207.5, 323, 275.5, 445.5, 416, 94.5, 478.5, 
    122.5, 107, 28.5, 274.5, 246.5, 456, 61.5, 104.5, 447.5, 25, 108.5, 189, 
    388, 255.5, 476, 196.5, 392, 172.5, 463, 455, 37, 356.5, 441.5, 300.5, 
    64.5, 264.5, 76, 10.5, 180.5, 171, 489, 303.5, 278.5, 17.5, 78.5, 25, 
    473.5, 140, 129.5, 421.5, 165, 238.5, 110.5, 53, 494, 87, 249.5, 386.5, 
    259.5, 213, 341.5, 297, 70, 283.5, 97.5, 134.5, 48, 174, 145, 229, 345, 
    134, 33, 123.5, 152, 111.5, 149, 126, 252, 279, 47.5, 417, 17.5, 158.5, 
    470.5, 12, 245.5, 220.5, 398.5, 5, 434, 240.5, 302.5, 4, 24, 400, 139, 
    72.5, 74, 284, 301.5, 419.5, 418.5, 335, 43.5, 71, 447, 192.5, 197, 199, 
    471.5, 245, 116.5, 489.5, 403.5, 87, 1.5, 149, 308, 400, 154.5, 242, 141, 
    457, 246, 165, 357, 385.5, 237.5, 431.5, 169.5, 39.5, 351.5, 88.5, 375, 
    395, 160, 322, 87.5, 357, 21, 59.5, 102, 138, 49, 6, 225.5, 51, 155, 
    33.5, 451.5, 310, 275.5, 92.5, 267, 22, 257.5, 124.5, 407.5, 495.5, 56.5, 
    77.5, 35, 408, 166.5, 410, 303, 326.5, 232.5, 391, 184, 254, 451, 286, 
    392, 0.5, 292.5, 117.5, 51.5, 448, 151.5, 3, 258, 427, 95.5, 25.5, 449.5, 
    353.5, 150, 357.5, 349, 207, 435.5, 384.5, 115.5, 102, 295, 419, 428.5, 
    27.5, 310, 113, 281.5, 261.5, 399, 174, 262, 192, 292, 314, 140, 443.5, 
    317, 398, 371, 413, 423.5, 320.5, 267, 74, 178, 116.5, 281.5, 113.5, 1, 
    397, 216, 296.5, 316, 145, 324, 126.5, 258, 106, 388, 157.5, 280.5, 150, 
    349.5, 72.5, 464.5, 489.5, 16, 281.5, 388, 387, 195, 311.5, 207.5, 462.5, 
    386, 386, 79, 167.5, 0, 80.5, 65, 216.5, 377, 381, 361.5, 201.5, 7.5, 
    120, 308, 396, 277.5, 88.5, 46.5, 127.5, 161, 11, 117, 177, 293, 5, 64.5, 
    488, 317, 272.5, 450.5, 203.5, 159, 29.5, 371, 159, 110, 436, 376, 487.5, 
    317.5, 237.5, 189, 325.5, 358, 497, 221.5, 135.5, 85.5, 268, 263.5, 
    246.5, 279, 380.5, 424, 72, 386, 488.5, 60.5, 203.5, 261, 11.5, 407, 420, 
    41, 278.5, 79.5, 151.5, 215, 456, 139.5, 33, 194, 328.5, 358.5, 52, 
    325.5, 80, 188, 411.5, 348, 451.5, 158.5, 127.5, 332.5, 83, 200, 219, 
    71.5, 260.5, 422.5, 333, 272, 330, 253.5, 313.5, 109, 333.5, 465.5, 
    324.5, 289.5, 105, 357.5, 483.5, 433.5, 216, 36, 259.5, 296, 224, 171, 
    144.5, 175.5, 330, 272, 8.5, 413, 472, 227.5, 484.5, 233, 150.5, 318, 5, 
    481, 72, 318.5, 90, 406, 284.5, 414.5, 196, 389.5, 272, 179.5, 323, 488, 
    216, 83, 284.5, 440, 254, 429, 116, 84, 201.5, 125, 497, 174, 352.5, 482, 
    407, 3.5, 300.5, 412.5, 484.5, 373, 231, 74.5, 279, 16, 489.5, 475, 
    405.5, 262, 155, 228.5, 250, 371, 312, 35, 311.5, 66, 464, 427.5, 150.5, 
    166, 52.5, 148, 340, 405.5, 130.5, 247.5, 409, 431.5, 160, 394, 304.5, 
    391.5, 468.5, 83.5, 407.5, 458.5, 58.5, 313, 220.5, 214, 42, 471, 85, 
    354, 6, 396.5, 420.5, 470.5, 324.5, 71.5, 136.5, 377.5, 219.5, 477, 
    283.5, 350.5, 224.5, 192.5, 282, 384.5, 86.5, 86.5, 276, 55.5, 170, 184, 
    14.5, 229, 497, 235, 443, 39, 206, 28.5, 393.5, 212.5, 425.5, 314, 183, 
    250.5, 385.5, 320, 128, 105.5, 297, 411.5, 456, 22, 104.5, 238, 406.5, 
    191.5, 324.5, 183, 247.5, 495, 367, 262, 224.5, 364, 497, 168, 403.5, 
    203.5, 196.5, 297.5, 416.5, 122.5, 111.5, 100, 373, 497.5, 420, 1, 103, 
    217.5, 413, 59, 239.5, 17.5, 297.5, 146.5, 209.5, 122, 329.5, 457, 117.5, 
    197, 219, 342, 61.5, 216.5, 10.5, 465, 420.5, 207.5, 262.5, 337, 330, 
    374.5, 437, 203, 372, 357.5, 204.5, 475.5, 75, 118, 35, 314.5, 136, 
    332.5, 461, 345.5, 455, 291, 302.5, 72.5, 488, 21.5, 415, 49.5, 238.5, 
    426, 15, 159, 133.5, 278, 496.5, 463.5, 153, 433.5, 167, 25, 291.5, 372, 
    1, 366.5, 490, 36, 181.5, 126, 369, 143, 472, 324, 434, 274.5, 397, 
    422.5, 296.5, 312.5, 472, 35.5, 238.5, 487.5, 194.5, 372, 265.5, 191, 
    336, 418.5, 125, 3.5, 444, 416.5, 375.5, 445.5, 283.5, 366, 481.5, 465, 
    492.5, 350.5, 108.5, 464.5, 175, 43, 239.5, 72.5, 465.5, 36.5, 385, 438, 
    72, 124, 425.5, 267, 496, 191.5, 458, 332.5, 110, 83.5, 336, 54.5, 0.5, 
    211.5, 0, 284, 77.5, 482, 249.5, 70.5, 333, 358, 35, 8, 401, 274.5, 81, 
    366.5, 311.5, 466, 305, 383.5, 90, 230.5, 150.5, 86.5, 422, 109, 419.5, 
    32.5, 193, 255.5, 87, 193.5, 467.5, 87.5, 477.5, 45.5, 69.5, 227.5, 116, 
    403, 86, 151, 411, 487, 426, 492.5, 354, 237.5, 458.5, 159, 121.5, 49, 
    390, 272.5, 136, 312, 381.5, 55.5, 344.5, 74.5, 311.5, 432, 268, 279, 
    19.5, 246, 324.5, 89.5, 474, 441, 492.5, 60, 92.5, 404, 47.5, 18.5, 
    396.5, 402, 256.5, 355.5, 61, 378.5, 404.5, 451.5, 151, 41, 263.5, 32.5, 
    97, 108.5, 107.5, 408.5, 40.5, 376, 188, 60.5, 122, 13, 150, 96.5, 454, 
    142.5, 156.5, 46.5, 46.5, 204, 65.5, 443, 106, 322, 299, 167.5, 201, 
    203.5, 119, 352, 245, 383, 384.5, 342, 491.5, 492, 250.5, 32.5, 368.5, 
    439, 93, 491, 452, 243.5, 87.5, 406, 386, 244, 452.5, 433, 448.5, 18.5, 
    376.5, 55, 341, 175.5, 223, 42, 379.5, 342, 394, 124.5, 225.5, 279, 
    466.5, 217, 271, 217.5, 250, 140, 156.5, 343, 131, 109, 87, 218.5, 15, 
    473, 463, 468, 406.5, 411.5, 486.5, 283, 467, 327.5, 459, 190, 370, 
    338.5, 32.5, 264, 463.5, 258, 43, 430.5, 475, 314.5, 148.5, 225.5, 454.5, 
    305, 69, 85.5, 414.5, 156, 304, 429.5, 129.5, 267, 398, 36, 179, 385, 
    319.5, 146.5, 212.5, 278.5, 336.5, 82.5, 117.5, 369, 347, 81.5, 127, 390, 
    12, 102.5, 204.5, 160.5, 328, 159.5, 466, 397, 245, 380.5, 53, 49.5, 
    310.5, 182.5, 317, 208.5, 219, 496.5, 93.5, 38.5, 143, 306.5, 317.5, 
    479.5, 389.5, 435.5, 348.5, 236.5, 17, 476, 126.5, 29, 78.5, 331.5, 
    189.5, 407, 491.5, 156, 304.5, 236.5, 36.5, 358, 286.5, 347, 41, 103.5, 
    55.5, 260, 100, 149.5, 299, 243.5, 456, 116.5, 223, 345.5, 52, 72, 82, 
    69, 48, 209, 98.5, 127, 41, 288.5, 34.5, 32.5, 444.5, 339, 269.5, 481, 
    197, 56, 328.5, 238, 160, 384.5, 498.5, 260, 34, 297.5, 3.5, 490, 414.5, 
    227, 336, 466.5, 299, 418.5, 36, 347.5, 128, 135, 475, 169, 423.5, 9.5, 
    202, 368, 348.5, 471.5, 349.5, 46, 28, 178, 284, 188, 63, 282.5, 448.5, 
    97, 80.5, 452.5, 87.5, 495, 180, 423.5, 462, 479.5, 342, 498, 327, 470.5, 
    133.5, 302.5, 139.5, 57, 312, 342, 425, 160.5, 313.5, 275, 206.5, 342, 
    453.5, 491, 30, 16.5, 274, 479, 113.5, 354.5, 432, 201.5, 349.5, 112, 
    125, 312, 91.5, 467.5, 310, 418.5, 438, 443.5, 221, 78, 1, 33.5, 420, 
    426.5, 194.5, 234, 201.5, 401.5, 76.5, 155, 392.5, 107, 172, 167, 86, 
    285.5, 21.5, 18, 487, 371.5, 130, 112.5, 183.5, 222, 80.5, 494, 140.5, 
    19, 438, 362, 97.5, 439, 396, 17.5, 365.5, 90.5, 252, 67.5, 492, 328.5, 
    223, 385, 435.5, 395, 52, 22, 181, 74, 40.5, 168.5, 445.5, 171, 281, 
    129.5, 393, 362, 124, 34, 381, 62, 396, 478.5, 1.5, 292.5, 496.5, 367.5, 
    383, 249, 435.5, 375, 78, 158.5, 260.5, 14, 54, 312.5, 36, 235, 386.5, 
    76.5, 403.5, 332.5, 248, 185, 462.5, 141, 47.5, 86.5, 175, 429, 149, 
    71.5, 408, 151, 364, 404.5, 19, 247, 154, 454.5, 122.5, 232, 113.5, 383, 
    246, 167.5, 196, 282, 402.5, 82.5, 359, 306.5, 415.5, 107, 491.5, 378.5, 
    248.5, 39.5, 465.5, 423.5, 468.5, 115, 495, 376.5, 266, 359, 281, 285, 
    106.5, 435, 240, 229, 167.5, 353.5, 112.5, 413.5, 21, 308.5, 196, 424, 
    391.5, 55.5, 230.5, 307.5, 163, 222.5, 186, 411.5, 262, 151.5, 335, 
    230.5, 266.5, 330.5, 107, 33, 189.5, 388.5, 318.5, 296.5, 324, 58.5, 
    25.5, 491.5, 412.5, 138.5, 405, 433.5, 447, 101.5, 357.5, 339, 157, 88.5, 
    146.5, 320.5, 311, 333, 232, 73, 484.5, 67.5, 303.5, 251.5, 398.5, 411, 
    284.5, 88, 299.5, 103.5, 385, 123.5, 162, 410.5, 115.5, 75, 49.5, 21, 
    8.5, 497, 122.5, 366.5, 336, 280, 455, 482.5, 100.5, 266.5, 315.5, 333, 
    339.5, 300.5, 401, 143.5, 52.5, 299.5, 55, 337, 388, 354.5, 441, 273, 
    478.5, 103, 184, 94, 178, 233.5, 115, 187, 230.5, 238, 54, 66.5, 18, 9.5, 
    49.5, 119, 276, 365.5, 452, 116, 166.5, 353.5, 260, 219, 153, 315, 56.5, 
    41, 170, 497.5, 314.5, 148.5, 101, 498.5, 242.5, 279.5, 232.5, 358, 467, 
    463, 96, 21, 30, 114.5, 31, 80, 233.5, 307, 446, 186, 423.5, 112.5, 39.5, 
    183.5, 332, 192.5, 499, 388.5, 234, 169, 386.5, 48.5, 317.5, 487.5, 47, 
    60.5, 267.5, 279.5, 419, 234.5, 243, 15, 255.5, 273, 129.5, 286.5, 353.5, 
    363.5, 94, 299.5, 49.5, 17.5, 412.5, 89, 201.5, 244.5, 281.5, 201, 133.5, 
    16, 370, 20, 64.5, 188, 8, 112, 249, 275.5, 392, 168, 10, 135, 183.5, 
    266, 408.5, 313, 52.5, 262, 176.5, 147, 62, 226.5, 165, 474.5, 315.5, 
    366.5, 219, 97.5, 68, 353, 113.5, 438, 373, 178, 126.5, 381, 290, 375.5, 
    157, 182.5, 44, 167, 317.5, 227.5, 433, 226.5, 41, 486, 488.5, 218, 133, 
    50.5, 444.5, 298, 25.5, 260, 165, 244.5, 358, 233, 98, 471.5, 171.5, 471, 
    150, 298.5, 352.5, 440.5, 174.5, 9.5, 123, 218.5, 177, 440.5, 446.5, 
    110.5, 167.5, 487.5, 96.5, 156, 205.5, 230, 207, 150.5, 28, 233, 411, 
    193.5, 478, 269, 427, 76, 240.5, 99, 47, 390.5, 398, 400, 331, 72.5, 410, 
    454, 291.5, 87, 395, 238, 197.5, 63, 225.5, 294.5, 219, 431.5, 24.5, 
    426.5, 82, 53, 159.5, 493, 246.5, 137.5, 262, 174, 214, 3, 273.5, 261, 
    393.5, 171.5, 161.5, 225, 244, 71.5, 179.5, 35.5, 159, 75, 273.5, 357, 
    138, 499, 151.5, 357.5, 431, 176.5, 284.5, 13, 229.5, 444.5, 6, 476.5, 
    82.5, 268.5, 150.5, 296.5, 271.5, 424.5, 58, 165.5, 96, 219.5, 391, 340, 
    291, 71, 375.5, 450.5, 146.5, 149.5, 307.5, 284.5, 149, 459.5, 142.5, 80, 
    136, 427.5, 93, 365.5, 372, 99.5, 342.5, 454.5, 368.5, 493.5, 251.5, 
    140.5, 418, 309.5, 306.5, 14, 29, 198, 354, 320.5, 269, 230, 271.5, 
    415.5, 379.5, 79, 200.5, 29, 38.5, 343.5, 109, 174.5, 271, 202.5, 40.5, 
    143, 302.5, 383, 98, 171.5, 376.5, 349.5, 312, 294.5, 159.5, 119, 309, 
    188.5, 317, 163, 9.5, 86.5, 393.5, 281, 2.5, 273.5, 360.5, 203, 302.5, 
    399, 47, 412, 74, 318, 115, 114.5, 461.5, 417.5, 498, 60, 89.5, 375, 410, 
    401.5, 170, 69.5, 21, 479, 258.5, 338, 142.5, 268, 424.5, 36, 49.5, 427, 
    310, 410, 130.5, 112.5, 309.5, 177.5, 25, 383.5, 496, 140, 498.5, 458, 
    58, 496.5, 18, 147.5, 372, 428, 49.5, 42, 497.5, 70.5, 21, 256, 408.5, 
    164, 24.5, 333.5, 200.5, 74, 261, 10.5, 484.5, 391.5, 123, 294, 69.5, 
    148.5, 177.5, 66, 288.5, 176, 24, 346.5, 173, 42.5, 494, 45.5, 470.5, 
    43.5, 87.5, 468.5, 114.5, 109, 225, 23.5, 273, 249.5, 357, 473.5, 324, 
    118, 484.5, 308.5, 10, 107.5, 102.5, 80, 256.5, 280.5, 146, 45, 457, 
    170.5, 392, 130.5, 213, 386, 176, 184, 430, 263.5, 152.5, 45, 373, 378, 
    68.5, 146.5, 128, 425.5, 120, 452, 44, 104.5, 261, 54.5, 212.5, 364, 
    134.5, 469.5, 144.5, 281, 14.5, 101.5, 451.5, 406.5, 232, 164.5, 293, 
    408.5, 349, 223.5, 172, 1.5, 268.5, 45.5, 380, 337, 192, 8, 263, 312.5, 
    460.5, 307.5, 417.5, 221.5, 362, 130.5, 86, 496.5, 100, 230.5, 278, 
    114.5, 332.5, 229.5, 21.5, 65, 394.5, 315, 473.5, 243.5, 38.5, 146, 
    245.5, 307.5, 191.5, 126, 145, 383.5, 134, 408.5, 196.5, 95, 216, 114, 
    317, 78, 244.5, 403, 75, 344.5, 133.5, 353, 459.5, 466, 83, 481.5, 31, 
    478, 296.5, 5, 222, 335.5, 151, 468, 143.5, 342.5, 94, 288.5, 226.5, 
    228.5, 197, 423, 323.5, 413, 37, 140.5, 491.5, 282, 43.5, 66.5, 127, 
    177.5, 420, 87, 144, 3, 68.5, 175.5, 481, 365.5, 180.5, 203.5, 201, 
    331.5, 171.5, 344.5, 174.5, 265.5, 133.5, 401, 494.5, 331, 324.5, 318, 
    244.5, 362, 459, 236, 144, 3, 303, 271.5, 180.5, 223, 358.5, 324.5, 
    226.5, 427, 0.5, 208, 292.5, 181, 411.5, 494, 12.5, 83, 339, 187, 349, 
    472.5, 88.5, 343.5, 304, 413, 162, 48.5, 275.5, 121, 285, 419.5, 124, 
    88.5, 191, 305, 311.5, 50, 129.5, 38.5, 477, 130, 246.5, 270, 311.5, 158, 
    264, 324.5, 241.5, 103, 12, 90.5, 76, 100.5, 434.5, 380, 14, 96.5, 429, 
    289.5, 217.5, 214.5, 209.5, 342, 303, 401, 147, 115, 451, 277, 153.5, 
    428.5, 407, 400.5, 198.5, 219, 59, 463, 43.5, 300.5, 66.5, 55.5, 391.5, 
    142.5, 156.5, 326, 23, 170.5, 423, 452.5, 460.5, 140.5, 167, 170, 482.5, 
    470, 71.5, 129.5, 85.5, 23, 406.5, 239.5, 451.5, 314, 140, 150.5, 33.5, 
    199, 113.5, 77, 0, 180, 132.5, 392, 323, 289, 218, 346, 460, 141.5, 
    298.5, 421, 282, 466, 91, 265, 436.5, 163, 395, 22, 186, 302, 261.5, 138, 
    116.5, 402, 288.5, 150, 101.5, 402.5, 227, 101.5, 83, 360, 493.5, 406, 
    149.5, 212, 252.5, 110, 353.5, 51.5, 31, 136, 17.5, 122, 401.5, 454, 
    285.5, 296.5, 476.5, 471.5, 98.5, 238.5, 109.5, 215, 140.5, 398.5, 365, 
    242.5, 301, 92.5, 344.5, 384, 453, 338, 290.5, 102.5, 50.5, 43, 212.5, 
    404.5, 95, 243.5, 41, 112.5, 366, 442.5, 67, 151.5, 239.5, 43.5, 123.5, 
    338.5, 282, 233.5, 54, 423, 132, 419.5, 165.5, 433.5, 12, 10, 317.5, 465, 
    348.5, 108.5, 68, 399.5, 152, 280.5, 304.5, 247, 24.5, 346, 360, 390.5, 
    289, 427, 42.5, 28.5, 471, 166.5, 367, 253.5, 400, 421, 176.5, 32, 340.5, 
    342.5, 465.5, 353, 353, 283.5, 318.5, 202, 392.5, 386.5, 102, 44.5, 167, 
    407, 292, 192, 253, 152, 82.5, 42, 79.5, 125.5, 71, 50.5, 292, 438.5, 
    304, 192, 360, 481, 224.5, 201, 324, 190.5, 54, 177.5, 474.5, 372.5, 380, 
    367.5, 259.5, 482, 412, 427, 389.5, 204.5, 119, 143, 357, 201.5, 185.5, 
    436.5, 327.5, 256.5, 487.5, 119.5, 195, 291.5, 312, 55.5, 273, 37, 256.5, 
    97, 227.5, 310.5, 274.5, 202.5, 183.5, 154.5, 70, 443, 137, 482.5, 370, 
    27, 187, 489, 170, 44.5, 191, 355.5, 481, 19, 112, 468.5, 138.5, 307.5, 
    260.5, 451, 363, 33.5, 488, 120, 131, 216, 430.5, 406, 418.5, 114.5, 61, 
    489, 58, 198, 471.5, 428.5, 225.5, 159, 418, 395.5, 204, 109.5, 251, 185, 
    128.5, 363.5, 154, 267.5, 171.5, 415, 218.5, 35, 448.5, 207, 155, 80, 
    423, 86, 486, 342, 200.5, 47, 331, 259, 245.5, 303, 187.5, 471, 462.5, 
    105.5, 366.5, 166.5, 215.5, 118, 352, 344, 481.5, 6.5, 111.5, 153, 421.5, 
    330.5, 188, 370.5, 37.5, 343.5, 450.5, 460.5, 429.5, 436.5, 302.5, 130.5, 
    483.5, 134, 389.5, 229.5, 437, 77.5, 200.5, 400, 183.5, 67, 66.5, 399, 
    185, 418.5, 243, 167, 425, 355, 320.5, 346.5, 185.5, 9, 217.5, 223, 
    352.5, 168, 184, 282, 105, 486.5, 413, 89, 121, 302.5, 318.5, 58.5, 380, 
    19, 458.5, 63.5, 86.5, 25, 462.5, 272, 444, 206, 439, 369, 61, 260, 216, 
    246.5, 269, 433.5, 470, 122, 102, 154, 404, 207, 141, 317.5, 296, 262, 
    120, 114.5, 320.5, 0.5, 134, 279, 64.5, 220.5, 304.5, 27, 492.5, 248.5, 
    233.5, 432, 117.5, 294.5, 192, 334, 41.5, 461.5, 268, 12, 83.5, 370.5, 
    166, 488, 77.5, 307, 305.5, 374, 69.5, 426, 489, 390, 426.5, 123, 169.5, 
    491, 344, 474, 18.5, 336.5, 222.5, 252, 269, 340.5, 47, 461.5, 175, 89, 
    423, 443.5, 101, 6.5, 314, 267.5, 494.5, 392, 75, 300.5, 266, 144.5, 
    226.5, 255.5, 35, 153, 378.5, 205, 144.5, 223, 179, 163, 60, 402, 415.5, 
    329, 243, 463, 290.5, 418.5, 52.5, 213.5, 362, 154, 220.5, 176, 421.5, 
    215.5, 68, 496.5, 16, 334.5, 141, 242.5, 90, 176.5, 396, 469, 381.5, 
    40.5, 192, 61, 204, 252, 463, 119.5, 81.5, 206.5, 83, 372, 125, 135.5, 
    86, 487, 289.5, 307, 163.5, 211.5, 22.5, 231.5, 208, 38.5, 66, 349.5, 
    281.5, 156, 26.5, 177.5, 125, 408, 218, 317, 469, 422, 69.5, 432.5, 42, 
    151, 139, 125.5, 23.5, 264.5, 261.5, 109.5, 252, 51.5, 416.5, 415.5, 263, 
    439.5, 147, 471.5, 478, 213.5, 321.5, 259.5, 370, 348, 437.5, 495, 256, 
    156, 312.5, 225.5, 78, 382.5, 158.5, 120.5, 33.5, 298, 246, 57, 62.5, 
    7.5, 167, 314.5, 59, 84, 230.5, 322.5, 23.5, 377.5, 294, 2, 91.5, 115.5, 
    262, 461.5, 464, 199.5, 457, 220, 355.5, 269.5, 446, 434, 152, 104.5, 55, 
    186, 402.5, 301, 243, 465.5, 309, 410.5, 280, 368.5, 494.5, 10.5, 191.5, 
    18.5, 388.5, 485.5, 20.5, 480.5, 101.5, 282.5, 442, 65.5, 482.5, 399, 
    286, 338, 169, 232.5, 272.5, 321, 337, 327.5, 7.5, 240, 129, 251, 205.5, 
    438.5, 161.5, 486, 307.5, 156.5, 497, 499, 175, 386, 484.5, 195.5, 366.5, 
    86.5, 478.5, 308.5, 152.5, 461, 208, 438.5, 299.5, 377, 171, 72.5, 198.5, 
    8.5, 400.5, 206, 248.5, 29.5, 457, 454.5, 468, 119, 440.5, 275.5, 275.5, 
    437.5, 275, 450.5, 323.5, 260, 146.5, 190.5, 346.5, 125.5, 499, 499, 87, 
    207.5, 438, 387, 84.5, 109.5, 459.5, 283.5, 118.5, 360, 490, 367.5, 390, 
    447.5, 322, 358.5, 66.5, 262.5, 134.5, 342.5, 200.5, 409.5, 293.5, 24.5, 
    169.5, 440.5, 215, 16.5, 66, 214.5, 15.5, 153.5, 422, 454, 40.5, 7, 64, 
    0.5, 290.5, 182.5, 361, 280.5, 50, 251, 228.5, 372.5, 110, 295, 135.5, 
    244.5, 138, 336, 154, 431.5, 360.5, 324, 372, 76, 340.5, 438, 290.5, 
    356.5, 92, 212.5, 310.5, 132.5, 219.5, 375, 133.5, 10.5, 58, 494.5, 
    291.5, 108.5, 246, 20, 481, 356, 315.5, 116.5, 101, 453.5, 453, 255.5, 
    385, 314, 79.5, 257.5, 390, 420, 196, 180.5, 276.5, 288, 393.5, 87.5, 
    420.5, 113.5, 463, 54, 124, 21, 49, 415.5, 129.5, 295, 436, 110.5, 151.5, 
    251.5, 227, 252.5, 205, 180.5, 8, 90.5, 494.5, 88, 348, 384.5, 8, 44.5, 
    65, 285, 332.5, 459, 373, 253, 72.5, 336, 307.5, 196.5, 357, 357, 112.5, 
    486.5, 152, 48.5, 97.5, 304, 300.5, 325, 57, 6, 5.5, 65, 97, 0, 153, 445, 
    384.5, 161.5, 489.5, 450, 446.5, 322.5, 409, 320, 76, 481.5, 156, 383.5, 
    178.5, 13, 241, 291.5, 0, 393, 340.5, 97.5, 197.5, 141, 422.5, 254.5, 
    147, 428, 320, 244, 428, 473, 189.5, 313, 135, 179.5, 263, 82, 2, 172.5, 
    402, 78.5, 154.5, 58, 462.5, 333.5, 71.5, 203.5, 125, 71.5, 97, 465.5, 
    169, 294.5, 106.5, 91.5, 49, 254, 19.5, 369, 498.5, 448, 342.5, 188.5, 
    261, 478, 368, 24, 60, 370.5, 197, 462.5, 449, 351.5, 20.5, 411.5, 185, 
    92, 115, 310.5, 164, 212.5, 276, 333, 7, 383, 424.5, 56.5, 137, 444.5, 
    426, 136, 392.5, 268.5, 324.5, 154, 247, 193, 178.5, 307, 63.5, 375.5, 
    269.5, 13, 227.5, 290.5, 425, 413, 383, 40.5, 223.5, 47, 253, 499.5, 380, 
    260.5, 382.5, 305, 317, 20, 250, 243, 156, 143, 12, 480.5, 297, 259, 
    173.5, 476, 66.5, 237.5, 351.5, 336, 251, 79, 127, 176, 492.5, 10, 217, 
    216, 57.5, 470.5, 215.5, 438, 231, 98.5, 243, 48, 118.5, 493.5, 291, 
    274.5, 136.5, 303.5, 255.5, 434, 62.5, 429, 410, 129, 167, 261.5, 465.5, 
    418, 341, 93, 94.5, 333.5, 103, 312, 50, 161, 282.5, 265.5, 99, 13.5, 
    364, 342.5, 62, 483, 336, 353.5, 257.5, 472.5, 157, 13, 407, 219.5, 
    442.5, 317, 349, 109.5, 79, 314.5, 28, 420.5, 407.5, 123, 254.5, 11, 435, 
    304.5, 172, 217.5, 70.5, 271, 231, 434.5, 113.5, 293.5, 417.5, 450, 147, 
    175.5, 423, 304, 189, 330, 23.5, 131.5, 147, 373, 241.5, 226, 187.5, 270, 
    147, 95.5, 393, 401.5, 106.5, 328, 206.5, 279, 45.5, 277, 50.5, 277, 
    211.5, 164.5, 70.5, 129.5, 114.5, 217.5, 305, 37.5, 22, 494, 368, 45.5, 
    126, 15, 419, 368, 241.5, 106.5, 138, 388.5, 202.5, 31, 290.5, 309.5, 
    359, 497, 88.5, 405, 274, 139.5, 182.5, 486, 304.5, 253.5, 115.5, 419.5, 
    471, 421, 457.5, 493, 415.5, 325.5, 39, 42, 340.5, 458.5, 410, 82.5, 65, 
    48, 471, 268, 79.5, 262, 77.5, 438.5, 259, 166.5, 344, 33.5, 306, 27, 
    19.5, 111, 280.5, 135.5, 30.5, 252, 57, 488, 245, 472.5, 313.5, 284.5, 
    14.5, 154.5, 243.5, 425, 237, 308.5, 473, 208, 76.5, 52.5, 470.5, 154.5, 
    491.5, 229.5, 321, 336, 263.5, 127.5, 363, 283, 238.5, 143.5, 419, 269, 
    395.5, 476, 257, 141, 449, 71, 426, 463.5, 225.5, 169.5, 388.5, 462.5, 
    478.5, 362, 171, 55.5, 415, 141.5, 210, 407, 371.5, 31, 243, 135, 158.5, 
    106, 418.5, 397.5, 250, 338, 166.5, 146, 314, 424, 287, 263, 495, 213.5, 
    227, 220.5, 383, 116, 183, 362, 478, 354.5, 417.5, 393.5, 496, 128, 
    300.5, 367.5, 159, 43.5, 3, 318, 150, 422, 215.5, 400.5, 260, 382.5, 
    46.5, 74, 306.5, 334, 337.5, 301.5, 47.5, 64.5, 22.5, 431, 180.5, 205.5, 
    293, 159, 60, 211, 53, 56.5, 339, 353.5, 424.5, 498.5, 397.5, 427.5, 317, 
    47.5, 349.5, 33, 448.5, 110, 415.5, 495, 184, 222.5, 329.5, 22, 24, 377, 
    86.5, 46.5, 308.5, 267.5, 252.5, 102, 427, 313, 313, 480, 369.5, 152.5, 
    334, 294, 151.5, 231.5, 222, 468.5, 279.5, 72, 1.5, 228, 182, 417.5, 
    223.5, 366.5, 140, 53, 388.5, 164.5, 430.5, 475.5, 211.5, 239, 243.5, 
    464, 341, 171, 277.5, 154.5, 151, 147, 307, 485, 441.5, 458.5, 217, 
    163.5, 427.5, 496.5, 236, 429.5, 224.5, 418, 347, 448, 285, 487.5, 1.5, 
    174, 152.5, 432, 149.5, 364, 171, 393, 328.5, 12.5, 64, 106, 167, 215.5, 
    253.5, 474.5, 201, 195, 433, 418, 359, 360.5, 414.5, 95.5, 290.5, 139.5, 
    14, 138, 88, 299, 125.5, 89.5, 473, 278.5, 21.5, 122.5, 142.5, 193, 16, 
    471.5, 205.5, 80.5, 78, 372.5, 296.5, 331.5, 347, 497.5, 27, 280.5, 416, 
    386.5, 141.5, 331, 482, 432, 470.5, 496, 70, 58.5, 295.5, 196, 148.5, 
    268.5, 474.5, 170, 391.5, 117.5, 363.5, 408, 89, 69, 489, 167, 442, 
    285.5, 499, 289.5, 283.5, 26.5, 70, 200, 413, 212, 31, 395.5, 144.5, 2, 
    391.5, 214.5, 61, 187.5, 411, 209.5, 456, 386, 380, 348, 3.5, 243.5, 
    256.5, 93, 312.5, 245.5, 260.5, 255, 31.5, 259.5, 44.5, 315.5, 286, 115, 
    15.5, 199.5, 327, 46.5, 95, 471.5, 49, 487, 186.5, 110, 174.5, 98, 319.5, 
    131, 484, 199.5, 479.5, 487.5, 443, 236, 81, 256, 481.5, 341.5, 11, 13.5, 
    101.5, 55.5, 329, 388, 171, 344.5, 88, 498, 391.5, 183, 470, 440.5, 
    170.5, 157, 50.5, 345, 255, 370, 476.5, 239, 70, 456, 227, 13, 192, 
    308.5, 269, 174, 150, 280, 187.5, 252, 336, 17, 140.5, 7, 361.5, 228.5, 
    5.5, 253.5, 412, 476, 194, 82.5, 133, 245, 428, 388.5, 115, 404.5, 128, 
    185, 360.5, 355, 198.5, 52.5, 163.5, 467.5, 227, 314, 248, 415, 66.5, 
    84.5, 432, 207, 92, 294, 435.5, 97.5, 47.5, 348, 73.5, 241.5, 430.5, 207, 
    486.5, 358.5, 95.5, 102, 263, 223.5, 287.5, 123.5, 79, 486, 176.5, 243, 
    454, 404, 57, 202.5, 319, 123.5, 287, 251.5, 331, 379, 45.5, 267, 477, 
    93, 115, 51, 335, 45.5, 258, 322, 404.5, 354, 424, 168, 78, 212, 292, 
    157, 198.5, 468.5, 400.5, 152.5, 373, 457.5, 355.5, 192, 81.5, 143, 
    443.5, 413, 22.5, 489.5, 180, 499.5, 82.5, 295, 50.5, 417.5, 341, 309, 
    240, 246, 163.5, 164, 414, 241.5, 376.5, 206, 399, 75, 175, 299.5, 228, 
    48, 257, 83.5, 240.5, 339, 226.5, 184.5, 252, 249.5, 174, 432.5, 249, 
    257, 227.5, 300, 175, 69, 109.5, 415, 315, 273, 79.5, 229, 14.5, 456, 
    435.5, 414, 31, 110.5, 213.5, 259, 159, 471, 343, 399.5, 310, 70, 84.5, 
    62.5, 319.5, 258.5, 495, 69, 15.5, 223, 369.5, 190.5, 292.5, 479.5, 106, 
    107.5, 252.5, 185.5, 337, 267.5, 141.5, 272.5, 181.5, 173, 383.5, 395.5, 
    432.5, 42.5, 366.5, 275.5, 442.5, 177, 346, 27, 239.5, 166, 285.5, 235, 
    235, 301.5, 458.5, 105, 492.5, 251, 84.5, 98.5, 359, 337.5, 284, 196.5, 
    105, 426, 469.5, 287, 99, 353, 182.5, 31.5, 396, 49, 307.5, 338.5, 226.5, 
    153.5, 365.5, 466.5, 319.5, 151, 201.5, 55, 453, 160.5, 160, 446, 411.5, 
    244.5, 44.5, 271, 82, 329, 467.5, 187.5, 255, 437, 474.5, 354, 290, 
    157.5, 386, 186, 207, 193.5, 24.5, 433.5, 347, 390, 400, 166.5, 41.5, 
    102, 221.5, 495, 262.5, 382, 441, 174.5, 126.5, 486, 445.5, 209, 315, 
    413, 396.5, 70.5, 350, 371.5, 425, 140.5, 29.5, 311, 327, 236.5, 4.5, 
    351.5, 170, 352, 242, 70.5, 19, 284, 172.5, 241, 279.5, 435.5, 123, 
    220.5, 110, 250, 206.5, 55.5, 459, 22, 469, 356, 92.5, 319, 228, 17.5, 
    460, 257.5, 329, 287, 494, 334, 139, 164.5, 186, 381.5, 235, 205, 165.5, 
    407.5, 446, 445.5, 343.5, 69.5, 166, 453.5, 319.5, 373, 9.5, 278.5, 
    395.5, 478.5, 135, 488.5, 298, 363, 6.5, 258, 120.5, 335.5, 45, 114.5, 
    169.5, 184, 279.5, 356, 65.5, 14.5, 61.5, 231.5, 422.5, 7.5, 177, 266, 
    77, 343.5, 219.5, 397, 217, 229, 175.5, 112.5, 208, 310.5, 101, 6, 174, 
    108, 264, 294.5, 443.5, 309, 409.5, 113.5, 493, 189, 469.5, 59, 203.5, 
    31, 290.5, 126.5, 39, 468, 392.5, 116.5, 311.5, 112, 13.5, 28.5, 341.5, 
    189.5, 141.5, 49.5, 0.5, 243, 55.5, 174.5, 351, 319.5, 469.5, 295, 129, 
    379.5, 408.5, 122.5, 68.5, 378.5, 181.5, 272.5, 410, 472.5, 399, 449.5, 
    440.5, 292, 66, 252.5, 404, 80, 281.5, 246, 270, 423, 296, 270.5, 166.5, 
    351.5, 445.5, 17.5, 171.5, 415.5, 313, 301, 295, 222, 423.5, 364, 100.5, 
    105.5, 137, 11, 78, 36.5, 460.5, 19, 328.5, 26.5, 271.5, 233, 107, 53, 
    479, 377, 476, 275, 148, 143, 127, 94, 161, 299, 9.5, 474, 100, 305, 196, 
    23.5, 169, 297, 129, 306, 308, 207.5, 343, 268.5, 226.5, 171.5, 295.5, 
    498, 404.5, 402.5, 51, 383.5, 280, 27.5, 159, 428.5, 170.5, 286.5, 23, 
    331.5, 85.5, 33, 306, 186, 338, 2, 209.5, 7.5, 299, 339, 314, 107, 46.5, 
    157, 375.5, 273, 328.5, 171, 271.5, 233, 74, 323, 117, 354.5, 350.5, 
    276.5, 283, 21.5, 63, 306.5, 353.5, 149, 339.5, 159.5, 335, 177.5, 161.5, 
    45, 185, 461, 384, 499.5, 68, 431, 156.5, 444, 204.5, 485, 115.5, 476, 
    218.5, 190, 299, 336, 44.5, 150, 112.5, 328, 171.5, 176, 134.5, 25.5, 
    325, 474, 185, 160.5, 152, 347, 205.5, 337.5, 308, 89.5, 337, 376.5, 21, 
    493.5, 321, 225.5, 479, 437, 202, 198, 127, 1, 34, 172, 151.5, 147, 0, 
    323.5, 323, 135, 349, 148.5, 109.5, 34.5, 309, 262, 381.5, 14.5, 99.5, 
    190, 104.5, 437, 67, 125.5, 430.5, 388.5, 351.5, 410, 325.5, 53.5, 108, 
    453, 54.5, 142.5, 125, 206.5, 289.5, 125.5, 30, 112.5, 261, 379, 261.5, 
    370.5, 414, 70.5, 132.5, 295.5, 85.5, 232.5, 486, 190.5, 169.5, 53, 316, 
    100.5, 442, 168, 11, 267.5, 221.5, 119, 220.5, 276.5, 262, 345.5, 483, 
    51.5, 471.5, 13.5, 164.5, 232.5, 393, 426, 103.5, 307, 497, 236, 102.5, 
    83, 469, 89, 273.5, 139, 142.5, 90, 239.5, 84.5, 258, 250.5, 352.5, 
    479.5, 370, 73, 256.5, 132, 419, 239.5, 184, 390.5, 253, 348.5, 123.5, 
    146, 274.5, 227, 453, 272, 463.5, 56, 355, 432.5, 145.5, 128.5, 71.5, 
    288, 218.5, 311.5, 373, 477, 62.5, 225.5, 457, 432.5, 299, 213.5, 65, 
    218, 453.5, 249, 109, 206.5, 97.5, 233, 353, 372.5, 460, 306.5, 145, 
    423.5, 363, 0, 356.5, 8.5, 129, 428.5, 297, 348, 240, 170, 325, 302.5, 
    396, 282, 235.5, 195, 496, 301, 413.5, 449.5, 50.5, 22.5, 156.5, 148.5, 
    255.5, 9.5, 21.5, 216, 316.5, 166.5, 139.5, 179.5, 167, 496.5, 188.5, 
    296, 425, 486, 144.5, 165.5, 156.5, 470, 468.5, 52.5, 252.5, 204, 247.5, 
    248.5, 5.5, 161.5, 198, 56, 184, 354.5, 204.5, 440, 364.5, 226, 156.5, 
    181, 393, 296.5, 361, 60, 293, 49.5, 356.5, 218, 36, 1.5, 383.5, 192.5, 
    471.5, 352, 245.5, 224, 56.5, 493, 473, 62.5, 155, 171, 119, 339.5, 26, 
    324, 280, 390.5, 50.5, 436.5, 72, 443.5, 233, 433, 4, 26, 483, 360.5, 
    244.5, 19, 362.5, 128.5, 211.5, 334, 481, 457.5, 58.5, 38, 451, 31.5, 
    100.5, 106, 202.5, 220, 445.5, 229, 44, 225.5, 119.5, 94.5, 162, 191.5, 
    38, 395, 125, 42.5, 421.5, 108, 403.5, 166.5, 127.5, 266, 295.5, 339.5, 
    100, 276.5, 297, 158.5, 315, 248, 190, 416, 354, 393, 136, 299.5, 122, 
    180, 25, 242, 275, 187.5, 434, 313, 82.5, 59, 356, 4.5, 167.5, 259.5, 
    171.5, 295, 25.5, 467, 134.5, 126, 244, 431.5, 285, 59, 179.5, 475, 475, 
    33.5, 368.5, 111.5, 333.5, 490.5, 291.5, 358.5, 233, 66.5, 46, 167, 380, 
    129, 226.5, 236.5, 134, 394, 496, 305.5, 189.5, 22, 273, 324, 148, 17, 
    256, 433, 76.5, 436, 408.5, 51.5, 470, 277, 163.5, 303.5, 268, 455, 
    162.5, 1.5, 22, 209, 168.5, 402.5, 338.5, 395.5, 139, 472.5, 290, 135.5, 
    278.5, 479.5, 157.5, 51.5, 304, 305.5, 69, 60, 239, 145.5, 496, 147.5, 
    197.5, 466, 425, 361, 270, 193.5, 316.5, 432.5, 195, 339, 141.5, 364, 
    241.5, 480, 259.5, 381, 453, 50, 16.5, 231.5, 29.5, 174, 283.5, 334, 480, 
    352.5, 394, 219.5, 498.5, 390.5, 367, 196.5, 357, 292.5, 57.5, 127, 486, 
    374.5, 60, 181.5, 213.5, 201.5, 45.5, 455.5, 182, 305.5, 336.5, 135, 
    355.5, 353, 367, 385.5, 27.5, 150.5, 219.5, 7.5, 3.5, 114, 227.5, 2.5, 5, 
    95, 199, 362.5, 387.5, 257, 490, 374, 131.5, 50, 55.5, 345.5, 252, 101.5, 
    301, 434.5, 407, 137.5, 69.5, 263, 491, 437, 149, 18.5, 88, 368.5, 26.5, 
    91.5, 483, 254, 94.5, 488.5, 349, 294, 351, 237, 51, 341.5, 111, 183, 
    391.5, 167, 28.5, 144, 268.5, 329.5, 78.5, 176, 467, 148.5, 439.5, 458.5, 
    85.5, 88.5, 477, 173.5, 457.5, 4, 265.5, 440.5, 258.5, 360.5, 429.5, 108, 
    154.5, 280.5, 345, 205.5, 122, 456.5, 388.5, 14, 124, 417, 158.5, 393, 
    246.5, 237, 69, 214, 385.5, 8.5, 172.5, 471.5, 97.5, 150, 145.5, 55, 
    154.5, 411, 496, 413.5, 271.5, 425.5, 21.5, 426, 206.5, 367, 132, 329, 
    324, 20.5, 343, 448, 438, 1.5, 341, 185, 239, 410.5, 399, 125, 419.5, 72, 
    96.5, 17, 222.5, 242, 72.5, 377.5, 153.5, 68.5, 291, 425.5, 494, 313, 
    352, 201, 180, 484, 30, 4.5, 5, 373.5, 453, 443, 375.5, 294, 128.5, 
    114.5, 205, 28, 239.5, 124.5, 100, 336.5, 142, 323, 79, 214.5, 200.5, 
    233, 283, 492, 158.5, 277.5, 305, 11, 479, 485.5, 495, 9, 490.5, 0.5, 
    382.5, 443.5, 443.5, 258, 238, 72.5, 373, 443, 100.5, 113, 67.5, 201, 
    449.5, 210, 24, 29, 424.5, 225, 262, 208, 217.5, 421, 485.5, 22.5, 432, 
    464.5, 8.5, 427.5, 474, 499, 428, 357, 443, 372, 115, 181, 444.5, 488, 
    124, 45, 101, 192, 246, 51, 402, 270.5, 80.5, 327, 496, 342.5, 35, 213.5, 
    264, 21, 236.5, 196.5, 486, 245, 124, 460, 244.5, 52, 317, 187.5, 424, 
    432.5, 369, 368.5, 421, 493, 414, 22.5, 185.5, 160.5, 73.5, 87.5, 431, 
    154, 414.5, 427, 497, 449.5, 141, 261.5, 471, 377.5, 458, 457, 123, 82, 
    417, 368, 134, 234.5, 56, 58.5, 167, 425, 427.5, 88, 418.5, 341.5, 110.5, 
    104, 2.5, 184.5, 191.5, 433.5, 339, 106.5, 361, 336.5, 56.5, 2.5, 98, 
    27.5, 380, 56, 484.5, 3.5, 138.5, 402, 371.5, 273, 136.5, 427.5, 331.5, 
    303.5, 353, 259.5, 391.5, 271.5, 101.5, 2.5, 375.5, 104, 187, 67.5, 38, 
    26.5, 174, 399, 363, 231, 401.5, 461, 258.5, 282, 17.5, 243.5, 285.5, 
    156, 145.5, 157.5, 429, 282.5, 85.5, 261, 86, 438.5, 21, 478, 210, 122.5, 
    481, 86, 226.5, 168, 153.5, 264.5, 195, 328, 164, 58, 59, 66, 19.5, 318, 
    348.5, 37, 62, 134, 193.5, 207.5, 292, 123, 490.5, 377.5, 384.5, 76.5, 
    316, 405.5, 55, 26.5, 28, 36, 113, 255, 204.5, 266.5, 20, 399.5, 95, 184, 
    457.5, 154.5, 250.5, 477.5, 472.5, 99, 14.5, 35, 233.5, 208.5, 242.5, 
    25.5, 331.5, 233.5, 403, 216, 310, 219.5, 121.5, 365.5, 246.5, 150, 
    401.5, 359.5, 405, 106, 126, 425, 6, 221.5, 109.5, 464, 376, 360.5, 
    441.5, 349, 460, 456.5, 384, 194, 165, 127, 219.5, 496.5, 360.5, 123, 
    213, 171, 342.5, 335, 36.5, 89, 485, 438, 448.5, 390.5, 44.5, 75, 316, 
    50.5, 297, 426, 14.5, 173, 286.5, 456.5, 22.5, 247, 413, 406.5, 441, 78, 
    33.5, 161, 75, 394.5, 284, 288, 65.5, 127, 123, 102, 216.5, 108.5, 40.5, 
    165, 499, 85, 240.5, 315.5, 136, 37.5, 241.5, 150.5, 211, 28.5, 107.5, 
    233.5, 275.5, 20.5, 140, 217, 99, 174, 378, 174, 69, 162, 462.5, 134.5, 
    289, 86, 237, 5.5, 194.5, 277.5, 171, 194, 362.5, 412, 9.5, 498.5, 450, 
    251, 149.5, 161, 279.5, 257.5, 394.5, 55.5, 278, 35, 272.5, 377.5, 209.5, 
    150.5, 51.5, 278.5, 313, 14.5, 413.5, 102, 100.5, 150.5, 108, 295, 428, 
    279.5, 489, 291, 191.5, 499, 290, 141.5, 250, 439.5, 302.5, 30, 197.5, 
    197.5, 86, 475.5, 233, 358.5, 353, 443, 9.5, 405, 221.5, 322.5, 419.5, 
    135.5, 425, 20, 286, 33.5, 315.5, 214.5, 313, 305, 5.5, 5, 304, 295.5, 
    146.5, 54.5, 235.5, 449.5, 85, 433, 147.5, 171, 409, 381, 30, 262.5, 324, 
    40, 167.5, 46, 362.5, 87.5, 181.5, 288, 108, 467.5, 322, 423.5, 182.5, 
    135, 229, 188, 140, 33.5, 484, 287, 88.5, 219.5, 237, 173.5, 153, 384.5, 
    345, 62, 265.5, 375, 324.5, 89.5, 415.5, 492.5, 136, 278.5, 80, 317.5, 
    66.5, 188, 285.5, 388.5, 112, 468, 24, 341, 156.5, 164.5, 375, 140.5, 
    452, 463.5, 360, 189, 137.5, 13.5, 73.5, 482.5, 75.5, 339.5, 358, 400.5, 
    429.5, 273.5, 393, 65.5, 52, 473, 383.5, 119, 161, 169, 8, 273.5, 137.5, 
    32.5, 114.5, 294, 197, 490, 434.5, 149.5, 453.5, 295, 338.5, 91.5, 308.5, 
    412.5, 74.5, 384.5, 252.5, 432.5, 285, 182, 206.5, 178, 248, 259, 151.5, 
    131.5, 378.5, 313, 300.5, 386.5, 86.5, 438, 419.5, 201.5, 232.5, 116.5, 
    191.5, 167, 266, 145.5, 462.5, 105, 237, 271, 17.5, 311.5, 156, 270, 
    244.5, 441, 452.5, 451.5, 119.5, 200.5, 211, 271.5, 332, 89.5, 84.5, 133, 
    476.5, 171.5, 71.5, 396, 373, 304, 13, 64.5, 471.5, 279.5, 210.5, 434, 
    384.5, 448, 205, 402.5, 259.5, 361.5, 173, 4.5, 302.5, 125.5, 456, 422.5, 
    326.5, 167, 194, 159, 257, 279, 292, 233.5, 450.5, 363.5, 129.5, 323.5, 
    168, 142.5, 388.5, 139.5, 422, 99, 73.5, 306.5, 47, 279, 209.5, 307, 
    140.5, 382.5, 312, 443.5, 8.5, 268, 366, 335, 435.5, 60.5, 494, 193, 
    339.5, 286.5, 426.5, 290, 150.5, 56, 114, 318.5, 199, 2.5, 458.5, 121, 
    102, 32, 428, 149.5, 311.5, 137.5, 456.5, 452, 20.5, 268.5, 395.5, 29.5, 
    37, 262, 364.5, 473, 323, 359, 166, 162.5, 146, 93, 453, 296.5, 149, 67, 
    115.5, 348, 69.5, 74, 469.5, 172, 106.5, 398, 321.5, 418, 36, 278.5, 
    370.5, 56.5, 47, 266.5, 86, 84.5, 29, 451, 57.5, 352, 310.5, 224, 14.5, 
    457, 317, 467.5, 254, 466.5, 35, 369.5, 315, 104.5, 444, 284.5, 277, 51, 
    183, 98.5, 469, 219, 377, 340, 276, 424.5, 106.5, 362.5, 9, 135.5, 313.5, 
    67, 487.5, 124.5, 291.5, 2.5, 82, 108.5, 470.5, 336, 75.5, 5.5, 206, 
    390.5, 110.5, 150.5, 175.5, 387.5, 201.5, 358.5, 486.5, 171, 77.5, 363.5, 
    11, 353.5, 288.5, 118, 216, 297.5, 253.5, 30, 365, 241.5, 155, 156.5, 
    244, 237, 265.5, 214.5, 73.5, 341, 220.5, 279.5, 232, 331, 430, 407.5, 
    218.5, 132, 266, 205, 303, 343.5, 69, 314.5, 197.5, 357.5, 432.5, 414, 
    155.5, 186.5, 444 ;
}
